module TriBitTest;

parameter Bits = 12;

logic Out[Bits - 1:0];
logic In[Bits -1 :0];

TriBitCheck TriBit(Out,In);





endmodule